library verilog;
use verilog.vl_types.all;
entity Pratica05_reg_1_bit_vlg_vec_tst is
end Pratica05_reg_1_bit_vlg_vec_tst;
