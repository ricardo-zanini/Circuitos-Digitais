library verilog;
use verilog.vl_types.all;
entity Pratica01 is
    port(
        co              : out    vl_logic;
        b               : in     vl_logic;
        a               : in     vl_logic;
        s               : out    vl_logic
    );
end Pratica01;
