library verilog;
use verilog.vl_types.all;
entity Pratica04_Adder_4bits_vlg_vec_tst is
end Pratica04_Adder_4bits_vlg_vec_tst;
