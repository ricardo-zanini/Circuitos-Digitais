library verilog;
use verilog.vl_types.all;
entity ProjetoFinalCD_vlg_vec_tst is
end ProjetoFinalCD_vlg_vec_tst;
