library verilog;
use verilog.vl_types.all;
entity Pratica06_cont_gen_1bit_vlg_check_tst is
    port(
        q               : in     vl_logic;
        sand            : in     vl_logic;
        sor             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Pratica06_cont_gen_1bit_vlg_check_tst;
