library verilog;
use verilog.vl_types.all;
entity Pratica01_vlg_vec_tst is
end Pratica01_vlg_vec_tst;
