library verilog;
use verilog.vl_types.all;
entity Pratica06_cont_gen_1bit_vlg_vec_tst is
end Pratica06_cont_gen_1bit_vlg_vec_tst;
