library verilog;
use verilog.vl_types.all;
entity Pratica04_Full_Adder_vlg_vec_tst is
end Pratica04_Full_Adder_vlg_vec_tst;
