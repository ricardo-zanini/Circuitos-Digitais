library verilog;
use verilog.vl_types.all;
entity Pratica06_cont_gen_4_bits_vlg_check_tst is
    port(
        q               : in     vl_logic_vector(0 to 3);
        sampler_rx      : in     vl_logic
    );
end Pratica06_cont_gen_4_bits_vlg_check_tst;
