library verilog;
use verilog.vl_types.all;
entity Pratica04_Bloco_Aritmetico_vlg_vec_tst is
end Pratica04_Bloco_Aritmetico_vlg_vec_tst;
