library verilog;
use verilog.vl_types.all;
entity Pratica05_div_freq_5_bits_vlg_vec_tst is
end Pratica05_div_freq_5_bits_vlg_vec_tst;
