library verilog;
use verilog.vl_types.all;
entity Pratica05_div_freq_1_bit is
    port(
        saida           : out    vl_logic;
        rst             : in     vl_logic;
        ck              : in     vl_logic
    );
end Pratica05_div_freq_1_bit;
