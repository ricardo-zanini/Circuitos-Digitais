library verilog;
use verilog.vl_types.all;
entity Pratica04_xor2_4bits_vlg_vec_tst is
end Pratica04_xor2_4bits_vlg_vec_tst;
