library verilog;
use verilog.vl_types.all;
entity Pratica05_reg_1_bit_vlg_check_tst is
    port(
        q               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Pratica05_reg_1_bit_vlg_check_tst;
